/*********************************** 
 * Show a Flying BOO on LCD.        *
 * Each image is 16x16 bits.        *
 ***********************************/

module lcd_control (LCD_CLK, RENDER_CLK, RENDER_DATA,
       LCD_DATA, LCD_ENABLE, LCD_RW, LCD_RSTN, LCD_CS1, LCD_CS2, LCD_DI);

	input  LCD_CLK;
    input  RENDER_CLK;
    input [0:15]  RENDER_DATA;
	output reg [7:0]  LCD_DATA;
	output LCD_ENABLE; 
	output reg LCD_RW;
	output LCD_RSTN;
	output reg LCD_CS1 = 1;
	output reg LCD_CS2 = 1;
	output reg LCD_DI;

	reg [7:0]  LCD_DATA_NEXT;
	reg LCD_RW_NEXT;
	reg LCD_DI_NEXT;
    reg LCD_CS1_NEXT, LCD_CS2_NEXT;
	
	reg [1:0]  STATE = Init, STATE_NEXT;
	reg [2:0]  X_PAGE, X_PAGE_NEXT;
	reg [5:0]  Y, Y_NEXT;
	reg [7:0]  PATTERN;
	reg [6:0]  INDEX, INDEX_NEXT; // extended
	
	reg START, START_NEXT;	
	reg NEW_PAGE, NEW_PAGE_NEXT;
	reg NEW_COL, NEW_COL_NEXT;
	reg [2:0] PAGE_COUNTER, PAGE_COUNTER_NEXT;
	reg [6:0] COL_COUNTER, COL_COUNTER_NEXT;
	reg ENABLE, ENABLE_NEXT;

	parameter Init = 2'd0, Set_StartLine = 2'd1, Clear_Screen = 2'd2, Copy_Image = 2'd3;
	
	assign LCD_ENABLE = LCD_CLK & ENABLE; // when ENABLE=1, LCD write can occur at falling edge of clock 
	assign LCD_RSTN = 1'b1;	
	
	always@(posedge LCD_CLK) begin
        STATE    <= STATE_NEXT;
        X_PAGE   <= X_PAGE_NEXT;
        Y  <= Y_NEXT;
        INDEX<= INDEX_NEXT;
        LCD_DI   <= LCD_DI_NEXT;
        LCD_RW   <= LCD_RW_NEXT;
        LCD_DATA <= LCD_DATA_NEXT;
        START <= START_NEXT;	
        NEW_PAGE <= NEW_PAGE_NEXT;
        NEW_COL <= NEW_COL_NEXT;
        COL_COUNTER <= COL_COUNTER_NEXT;
        PAGE_COUNTER <= PAGE_COUNTER_NEXT;
        ENABLE <= ENABLE_NEXT;
        LCD_CS1 <= LCD_CS1_NEXT;
        LCD_CS2 <= LCD_CS2_NEXT;
	end

	always @(*) begin
		// default assignments
		STATE_NEXT  = STATE;
		X_PAGE_NEXT = X_PAGE;
		Y_NEXT = Y;
		INDEX_NEXT = INDEX;
		LCD_DI_NEXT = LCD_DI;
		LCD_RW_NEXT = LCD_RW;
		LCD_DATA_NEXT = LCD_DATA;	
		COL_COUNTER_NEXT = COL_COUNTER; 
		PAGE_COUNTER_NEXT = PAGE_COUNTER;
        LCD_CS1_NEXT = LCD_CS1;
        LCD_CS2_NEXT = LCD_CS2;
		START_NEXT =	1'b0;	
		NEW_PAGE_NEXT = 1'b0;
		NEW_COL_NEXT = 1'b0;	
		ENABLE_NEXT = 1'b0;
        
		case(STATE)
			Init: begin  //initial state
				STATE_NEXT =  Set_StartLine;
				// prepare LCD instruction to turn display on
				LCD_DI_NEXT = 1'b0;
				LCD_RW_NEXT = 1'b0;
				LCD_DATA_NEXT = 8'b0011111_1;
				ENABLE_NEXT = 1'b1;
			end
			Set_StartLine: begin //set start line
				STATE_NEXT = Clear_Screen;
				// prepare LCD instruction to set start line
				LCD_DI_NEXT = 1'b0;
				LCD_RW_NEXT = 1'b0;
				LCD_DATA_NEXT = 8'b11_000000; // start line = 0
				ENABLE_NEXT = 1'b1;
				START_NEXT = 1'b1;
			end
			Clear_Screen: begin
				if (START) begin
					NEW_PAGE_NEXT = 1'b1;
					PAGE_COUNTER_NEXT = 0;
					COL_COUNTER_NEXT = 0;
					X_PAGE_NEXT = 0; // set initial X address
					Y_NEXT = 0; // set initial Y address
				end else	
				if (NEW_PAGE) begin
					// prepare LCD instruction to move to new page
					LCD_DI_NEXT = 1'b0;
					LCD_RW_NEXT = 1'd0;
					LCD_DATA_NEXT = {5'b10111, X_PAGE};
					ENABLE_NEXT = 1'b1;
					NEW_COL_NEXT = 1'b1;
				end else if (NEW_COL) begin 
					// prepare LCD instruction to move to column 0 
					LCD_DI_NEXT    = 1'b0;
					LCD_RW_NEXT    = 1'd0;
					LCD_DATA_NEXT  = 8'b01_000000; // to move to column 0
					ENABLE_NEXT = 1'b1;
				end else if (COL_COUNTER < 64) begin
					// prepare LCD instruction to write 00000000 into display RAM
					LCD_DI_NEXT    = 1'b1;
					LCD_RW_NEXT    = 1'd0;
					LCD_DATA_NEXT  = 8'b00000000;
					ENABLE_NEXT = 1'b1;
					COL_COUNTER_NEXT = COL_COUNTER + 1;
				end else begin
					if (PAGE_COUNTER == 7) begin // last page of screen
						STATE_NEXT = Copy_Image;
						START_NEXT = 1'b1;
					end else begin
						// prepare to change page
						X_PAGE_NEXT  = X_PAGE + 1;
						NEW_PAGE_NEXT = 1'b1;
						PAGE_COUNTER_NEXT = PAGE_COUNTER + 1;
						COL_COUNTER_NEXT = 0;
					end
				end
			end						
			Copy_Image: begin // write image pattern into LCD RAM
				if (START) begin
					NEW_PAGE_NEXT = 1'b1;
					X_PAGE_NEXT = 0;  // image initial X address
					Y_NEXT = 0; // image initial Y address
					PAGE_COUNTER_NEXT = 0;
					COL_COUNTER_NEXT = 0;
                    INDEX_NEXT = 0; // pattern initial index
                    // Draw left side of the LCD
                    LCD_CS1_NEXT = 1'b1;
                    LCD_CS2_NEXT = 1'b0;
				end else if (NEW_PAGE) begin
					// prepare LCD instruction to move to new page 
					LCD_DI_NEXT = 1'b0;
					LCD_RW_NEXT = 1'b0;
					LCD_DATA_NEXT = {5'b10111, X_PAGE}; 
					ENABLE_NEXT = 1'b1;
					NEW_COL_NEXT = 1'b1;
				end else if (NEW_COL) begin
					// prepare LCD instruction to move to new column
					LCD_DI_NEXT = 1'b0;
					LCD_RW_NEXT = 1'b0;
					LCD_DATA_NEXT = {2'b01,Y};
					ENABLE_NEXT = 1'b1;
				end else if (COL_COUNTER < 64) begin //load image 1 byte at a time, 16 is the width of image
					// prepare LCD instruction to write image data into display RAM
					LCD_DI_NEXT = 1'b1;
					LCD_RW_NEXT = 1'b0;
					LCD_DATA_NEXT = PATTERN;
					ENABLE_NEXT = 1'b1;
					INDEX_NEXT = INDEX + 1;
					COL_COUNTER_NEXT = COL_COUNTER + 1;
				end else begin
                    if (LCD_CS1) begin
                        // change to right side of LCD
                        LCD_CS1_NEXT = 1'b0;
                        LCD_CS2_NEXT = 1'b1;
                        COL_COUNTER_NEXT = 0;
                        NEW_PAGE_NEXT = 1'b1;
                    end
					else if (PAGE_COUNTER == 7) begin // last page of image
						START_NEXT = 1'b1;
					end else begin
						// prepare to change page
						X_PAGE_NEXT = X_PAGE + 1;
						NEW_PAGE_NEXT = 1'b1;
						PAGE_COUNTER_NEXT = PAGE_COUNTER + 1;
						COL_COUNTER_NEXT = 0;
                        LCD_CS1_NEXT = 1'b1;
                        LCD_CS2_NEXT = 1'b0;
					end
				end				
			end
			default: STATE_NEXT = Init;
		endcase
    end
    
    parameter AIR = 4'b0000,
              WALL = 4'b0001,
              STONE = 4'b0010,
              BOMB = 4'b1111,
              BOMB_EXPLODE = 4'b1000;
    
    reg [0:159]  MAP, MAP_NEXT;
    reg [0:5]   GSTATE = 0, GSTATE_NEXT;
    reg [11:0]  P1_POS, P2_POS;
    reg [11:0]  P1_POS_NEXT, P2_POS_NEXT;
    reg [1:0]   P1_DIR, P2_DIR, P1_DIR_NEXT, P2_DIR_NEXT;
    
    always @(posedge RENDER_CLK) begin
        MAP <= MAP_NEXT;
        GSTATE <= GSTATE_NEXT;
        P1_POS <= P1_POS_NEXT;
        P2_POS <= P2_POS_NEXT;
        P1_DIR <= P1_DIR_NEXT;
        P2_DIR <= P2_DIR_NEXT;
    end
    
    
    
    reg [2:0]  TX, TY; // Tile position
    reg [3:0]  IX, IY; // Image index
    reg [5:0]  PX; // Pixel X
    reg [3:0]  IMAGE;
    reg [0:143]  IMG_OUT;
    integer i;
    integer PL_X, PL_Y;
    integer OF_X, OF_Y;
    
    always @(*) begin
        IMAGE = 0;
            
        for (i = 7; i >= 0; i = i - 1) begin
            PX = X_PAGE * 8 + i;
            
            if (PX == 0 || PX == 63 || INDEX == 0 || INDEX == 127 || INDEX == 99) begin
                PATTERN[i] = 1'b1; // Black outter frame
            end
            else if (PX == 1 || PX == 62 || INDEX == 1 || INDEX == 126 || INDEX == 98 || INDEX == 100) begin
                PATTERN[i] = 1'b0; // White margin
            end
            else if (INDEX > 100) begin
                if (PX < 8 || PX >= 56) PATTERN[i] = 1'b0;
                else begin
                    case (GSTATE[0:1])
                        2'b00: begin
                            PATTERN[i] = PRESS_ZERO_TO_START[(PX-8) * 25 + (INDEX - 101)];
                        end
                        
                        2'b01: begin
                            case (GSTATE[2:3])
                                2'b00: PATTERN[i] = BATTLE[(PX-8) * 25 + (INDEX - 101)];
                                2'b01: begin
                                    if (PX[5] == 1'b0)
                                        PATTERN[i] = CD_1[(PX-8) * 25 + (INDEX - 101)];
                                    else
                                        PATTERN[i] = SEC_TO_START[(PX-32) * 25 + (INDEX - 101)];
                                end
                                2'b10: begin
                                    if (PX[5] == 1'b0)
                                        PATTERN[i] = CD_2[(PX-8) * 25 + (INDEX - 101)];
                                    else
                                        PATTERN[i] = SEC_TO_START[(PX-32) * 25 + (INDEX - 101)];
                                end
                                2'b11: begin
                                    if (PX[5] == 1'b0)
                                        PATTERN[i] = CD_3[(PX-8) * 25 + (INDEX - 101)];
                                    else
                                        PATTERN[i] = SEC_TO_START[(PX-32) * 25 + (INDEX - 101)];
                                end
                            endcase
                        end
                        
                        2'b10: begin
                            PATTERN[i] = GUIDE[(PX-8) * 25 + (INDEX - 101)];
                        end
                        
                        2'b11: begin
                            if (GSTATE[4:5] == 2'b10)
                                PATTERN[i] = WIN[(PX-8) * 25 + (INDEX - 101)];
                            else
                                PATTERN[i] = LOSE[(PX-8) * 25 + (INDEX - 101)];
                        end
                    endcase
                end
            end
            else begin
                // Main game map
                TX = (PX - 2) / 12;
                TY = (INDEX - 2) / 12;
                IX = (PX - 2) % 12;
                IY = (INDEX - 2) % 12;
                
                IMAGE = MAP[{TX, TY, 2'b00} +: 4];
                
                IMG_OUT = 0;
                if (IMAGE == WALL)
                    IMG_OUT = {12'b111111111111,
                               12'b100001000001,
                               12'b111111111111,
                               12'b100010001001,
                               12'b111111111111,
                               12'b101000010001,
                               12'b101000010001,
                               12'b111111111111,
                               12'b100010000101,
                               12'b111111111111,
                               12'b101000010001,
                               12'b111111111111};
                
                else if (IMAGE == STONE)
                    IMG_OUT = {12'b111111111111,
                               12'b100000000001,
                               12'b101111111101,
                               12'b101000000101,
                               12'b101000000101,
                               12'b101000000101,
                               12'b101000000101,
                               12'b101000000101,
                               12'b101000000101,
                               12'b101111111101,
                               12'b100000000001,
                               12'b111111111111};
                
                else if (IMAGE[3]) begin
                    if (IMAGE[0])
                        IMG_OUT = {12'b000000000110,
                                   12'b000000001001,
                                   12'b000111110001,
                                   12'b001001111000,
                                   12'b010000111000,
                                   12'b100000011100,
                                   12'b100000001100,
                                   12'b100000000100,
                                   12'b010000000100,
                                   12'b010000001000,
                                   12'b001000010000,
                                   12'b000111100000};
                    
                    else if (IMAGE[2:0] != 0)
                        IMG_OUT = {12'b000000000000,
                                   12'b000000000100,
                                   12'b000000001010,
                                   12'b000111110010,
                                   12'b001001110000,
                                   12'b010000110000,
                                   12'b010000011000,
                                   12'b010000001000,
                                   12'b010000001000,
                                   12'b001000010000,
                                   12'b000111100000,
                                   12'b000000000000};
                    
                    else
                        IMG_OUT = {12'b001010011010,
                                   12'b010100101010,
                                   12'b000111010011,
                                   12'b001001010101,
                                   12'b100110010010,
                                   12'b000111001010,
                                   12'b010101100111,
                                   12'b101101010111,
                                   12'b001011100101,
                                   12'b010010100101,
                                   12'b010100100100,
                                   12'b010010100101};
                end
                
                PATTERN[i] = IMG_OUT[12*IX + IY];
                
                
                // Player 1
                case (P1_DIR)
                        2'b00:
                            IMG_OUT = {12'b001111111100,
                                       12'b010000000010,
                                       12'b010000000010,
                                       12'b010000000010,
                                       12'b010000000010,
                                       12'b010000000010,
                                       12'b110000000011,
                                       12'b010000000010,
                                       12'b001111111100,
                                       12'b001010010100,
                                       12'b010010010010,
                                       12'b001100001100};
                        2'b01:
                            IMG_OUT = {12'b001111111100,
                                       12'b010000000010,
                                       12'b010000000010,
                                       12'b010010010010,
                                       12'b010010010010,
                                       12'b010010010010,
                                       12'b110000000011,
                                       12'b010000000010,
                                       12'b001111111100,
                                       12'b001010010100,
                                       12'b010010010010,
                                       12'b001100001100};
                        2'b10:
                            IMG_OUT = {12'b000111111000,
                                       12'b001000000100,
                                       12'b001000000100,
                                       12'b001010000100,
                                       12'b001010000100,
                                       12'b001010000100,
                                       12'b001000000100,
                                       12'b001000000100,
                                       12'b000111111000,
                                       12'b000001010000,
                                       12'b000010010000,
                                       12'b000001100000};
                        2'b11:
                            IMG_OUT = {12'b000111111000,
                                       12'b001000000100,
                                       12'b001000000100,
                                       12'b001000010100,
                                       12'b001000010100,
                                       12'b001000010100,
                                       12'b001000000100,
                                       12'b001000000100,
                                       12'b000111111000,
                                       12'b000010100000,
                                       12'b000010010000,
                                       12'b000001100000};
                    endcase
                
                PL_X = P1_POS[11:9] * 12 + P1_POS[8:6] * 2 + 2;
                PL_Y = P1_POS[5:3] * 12 + P1_POS[2:0] * 2 + 2;
                OF_X = PX - PL_X;
                OF_Y = INDEX - PL_Y;
                
                if (OF_X >= 0 && OF_X < 12 && OF_Y >= 0 && OF_Y < 12)
                    PATTERN[i] = IMG_OUT[OF_X * 12 + OF_Y];
                          
                     
                     //  player 2
                     
                     case (P2_DIR)
                        2'b00:
                            IMG_OUT = {12'b001111111100,
                                       12'b011111111110,
                                       12'b011111111110,
                                       12'b010000000010,
                                       12'b010000000010,
                                       12'b010000000010,
                                       12'b110000000011,
                                       12'b010000000010,
                                       12'b001111111100,
                                       12'b001010010100,
                                       12'b010010010010,
                                       12'b001100001100};
                        2'b01:
                            IMG_OUT = {12'b001111111100,
                                       12'b011111111110,
                                       12'b011111111110,
                                       12'b010000000010,
                                       12'b010010010010,
                                       12'b010010010010,
                                       12'b110010010011,
                                       12'b010000000010,
                                       12'b001111111100,
                                       12'b001010010100,
                                       12'b010010010010,
                                       12'b001100001100};
                        2'b10:
                            IMG_OUT = {12'b000111111000,
                                       12'b001111111100,
                                       12'b001111111100,
                                       12'b001000000100,
                                       12'b001010000100,
                                       12'b001010000100,
                                       12'b001010000100,
                                       12'b001000000100,
                                       12'b000111111000,
                                       12'b000001010000,
                                       12'b000010010000,
                                       12'b000001100000};
                        2'b11:
                            IMG_OUT = {12'b000111111000,
                                       12'b001111111100,
                                       12'b001111111100,
                                       12'b001000000100,
                                       12'b001000010100,
                                       12'b001000010100,
                                       12'b001000010100,
                                       12'b001000000100,
                                       12'b000111111000,
                                       12'b000010100000,
                                       12'b000010010000,
                                       12'b000001100000};
                    endcase
                
                PL_X = P2_POS[11:9] * 12 + P2_POS[8:6] * 2 + 2;
                PL_Y = P2_POS[5:3] * 12 + P2_POS[2:0] * 2 + 2;
                OF_X = PX - PL_X;
                OF_Y = INDEX - PL_Y;
                
                if (OF_X >= 0 && OF_X < 12 && OF_Y >= 0 && OF_Y < 12)
                    PATTERN[i] = IMG_OUT[OF_X * 12 + OF_Y];
                     
                     
            end
        end
    end
    
    always @(*) begin
        MAP_NEXT = MAP;
        GSTATE_NEXT = GSTATE;
        P1_POS_NEXT = P1_POS;
        P2_POS_NEXT = P2_POS;
        P1_DIR_NEXT = P1_DIR;
        P2_DIR_NEXT = P2_DIR;
        
        if (RENDER_DATA[0]) begin
            case (RENDER_DATA[1:2])
                2'b00: begin
                    MAP_NEXT[RENDER_DATA[3:8] * 4 +: 4] = RENDER_DATA[9:12];
                end
                
                2'b01: begin
                
                end
                
                2'b10: begin
                    GSTATE_NEXT = RENDER_DATA[3:8];
                end
                
                2'b11: begin
                
                end
            endcase
        end
        else begin
            if (RENDER_DATA[13] == 1'b0) begin
                P1_POS_NEXT = RENDER_DATA[1:12];
                P1_DIR_NEXT = RENDER_DATA[14:15];
            end
            else begin
                P2_POS_NEXT = RENDER_DATA[1:12];
                P2_DIR_NEXT = RENDER_DATA[14:15];
            end
        end
    end
    
    wire [0:599] CD_3 // 25 x 24
        = {25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000011111100000000000,
           25'b0000000111111110000000000,
           25'b0000000110001111000000000,
           25'b0000000000000111000000000,
           25'b0000000000000111000000000,
           25'b0000000000000111000000000,
           25'b0000000000001110000000000,
           25'b0000000011111100000000000,
           25'b0000000011111110000000000,
           25'b0000000000001111000000000,
           25'b0000000000000111000000000,
           25'b0000000000000111000000000,
           25'b0000000000000111000000000,
           25'b0000001100001111000000000,
           25'b0000001111111110000000000,
           25'b0000000111111100000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000};
    
    wire [0:599] CD_2
        = {25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000111110000000000,
           25'b0000000011111111000000000,
           25'b0000000111000011100000000,
           25'b0000000110000001100000000,
           25'b0000000000000001100000000,
           25'b0000000000000011100000000,
           25'b0000000000000111000000000,
           25'b0000000000001110000000000,
           25'b0000000000011100000000000,
           25'b0000000000111000000000000,
           25'b0000000001110000000000000,
           25'b0000000011100000000000000,
           25'b0000000111111111100000000,
           25'b0000000111111111100000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000};
           
    wire [0:599] CD_1
        = {25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000111000000000000,
           25'b0000000111111000000000000,
           25'b0000000110111000000000000,
           25'b0000000000111000000000000,
           25'b0000000000111000000000000,
           25'b0000000000111000000000000,
           25'b0000000000111000000000000,
           25'b0000000000111000000000000,
           25'b0000000000111000000000000,
           25'b0000000000111000000000000,
           25'b0000000000111000000000000,
           25'b0000000000111000000000000,
           25'b0000000111111111000000000,
           25'b0000000111111111000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000};
           
    wire [0:599] SEC_TO_START
        = {25'b0000000000000000000000000,
           25'b0000111100111110011111000,
           25'b0001000000100000100000000,
           25'b0000111100111110100000000,
           25'b0000000010100000100000000,
           25'b0001111100111110011111000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000111110111100000000,
           25'b0000000001000100100000000,
           25'b0000000001000100100000000,
           25'b0000000001000100100000000,
           25'b0000000001000111100000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0011101111101100111011111,
           25'b0100000010010010100100100,
           25'b0011100010011110111000100,
           25'b0000010010010010101000100,
           25'b0111100010010010100100100,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000};
           
    wire [0:1199] BATTLE
        = {25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b1110001100111011101000111,
           25'b1001010010010001001000100,
           25'b1110010010010001001000111,
           25'b1001011110010001001000100,
           25'b1001010010010001001000100,
           25'b1110010010010001001110111,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000001000100000000000,
           25'b0000000001000100000000000,
           25'b0000000001000100000000000,
           25'b0000000001000100000000000,
           25'b0000000001000100000000000,
           25'b0000000000000000000000000,
           25'b0000000001000100000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000};
           
    wire [0:1199] GUIDE
        = {25'b0000000000000011111110000,
           25'b0000010000000100000001000,
           25'b0000111000000101111101000,
           25'b0001010100000101000001000,
           25'b0000010000000101111101000,
           25'b0000010000000101000101000,
           25'b0000010000000101111101000,
           25'b0000010000000100000001000,
           25'b0000010000000011111110000,
           25'b0000000000000000000000000,
           25'b0000000000000011111110000,
           25'b0000010000000100000001000,
           25'b0000010000000101111101000,
           25'b0000010000000101000001000,
           25'b0000010000000101111101000,
           25'b0001010100000100000101000,
           25'b0000111000000101111101000,
           25'b0000010000000100000001000,
           25'b0000000000000011111110000,
           25'b0000000000000000000000000,
           25'b0000000000000011111110000,
           25'b0000000000000100000001000,
           25'b0000100000000101111101000,
           25'b0001000000000100000101000,
           25'b0011111110000101111101000,
           25'b0001000000000101000001000,
           25'b0000100000000101111101000,
           25'b0000000000000100000001000,
           25'b0000000000000011111110000,
           25'b0000000000000000000000000,
           25'b0000000000000011111110000,
           25'b0000000000000100000001000,
           25'b0000001000000101111101000,
           25'b0000000100000101000101000,
           25'b0011111110000101111101000,
           25'b0000000100000101000101000,
           25'b0000001000000101111101000,
           25'b0000000000000100000001000,
           25'b0000000000000011111110000,
           25'b0000000000000000000000000,
           25'b0000000011000011111110000,
           25'b0001111100100100000001000,
           25'b0010011100000100111001000,
           25'b0100001110000101000101000,
           25'b0100000110000101000101000,
           25'b0100000010000100111001000,
           25'b0010000100000100000001000,
           25'b0001111000000011111110000};
    
    wire [0:1199] PRESS_ZERO_TO_START
        = {25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0111101110011101111011110,
           25'b0100101001010001000010000,
           25'b0111101110011101111011110,
           25'b0100001010010000001000010,
           25'b0100001001011101111011110,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000011111111100000000,
           25'b0000000100000000010000000,
           25'b0000000100011100010000000,
           25'b0000000100100010010000000,
           25'b0000000100100010010000000,
           25'b0000000100100010010000000,
           25'b0000000100100010010000000,
           25'b0000000100011100010000000,
           25'b0000000100000000010000000,
           25'b0000000011111111100000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000111111100000000000,
           25'b0000000000100000000000000,
           25'b0000000000100011110000000,
           25'b0000000000100010010000000,
           25'b0000000000100010010000000,
           25'b0000000000100011110000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0011101111101100111011111,
           25'b0100000010010010100100100,
           25'b0011100010011110111000100,
           25'b0000010010010010100100100,
           25'b0111100010010010100010100,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000};
    
    wire [0:1199] WIN
        = {25'b0010001001111100100001000,
           25'b0010001010000010100001000,
           25'b0001010010000010100001000,
           25'b0001010010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100001111100011110000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0100100101111101100001000,
           25'b0100100100010001010001000,
           25'b0100100100010001010001000,
           25'b0010101000010001001001000,
           25'b0010101000010001001001000,
           25'b0010101000010001000101000,
           25'b0010101000010001000101000,
           25'b0001010001111101000011000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000101111111111111010000,
           25'b0001011000000000001101000,
           25'b0001001000000000001001000,
           25'b0001001100000000011001000,
           25'b0000110100000000010110000,
           25'b0000000100000000010000000,
           25'b0000000010000000100000000,
           25'b0000000001000001000000000,
           25'b0000000000111110000000000,
           25'b0000000000010100000000000,
           25'b0000000000010100000000000,
           25'b0000000000010100000000000,
           25'b0000000000010100000000000,
           25'b0000000000100010000000000,
           25'b0000001111111111111000000,
           25'b0000001000000000001000000,
           25'b0000001111111111111000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000};
           
    wire [0:1199] LOSE
        = {25'b0010001001111100100001000,
           25'b0010001010000010100001000,
           25'b0001010010000010100001000,
           25'b0001010010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100010000010100001000,
           25'b0000100001111100011110000,
           25'b0000000000000000000000000,
           25'b1000000111100011110011111,
           25'b1000001000010100000010000,
           25'b1000001000010100000010000,
           25'b1000001000010100000010000,
           25'b1000001000010011100011110,
           25'b1000001000010000010010000,
           25'b1000001000010000010010000,
           25'b1000001000010000010010000,
           25'b1000001000010000010010000,
           25'b1111100111100111100011111,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000000000000000000,
           25'b0000000000111100000000000,
           25'b0000000001000010000000000,
           25'b0000000000111100000000000,
           25'b0000000000000000000000000,
           25'b0000000000111110000000000,
           25'b0000000011000001000000000,
           25'b0001100100000000100110000,
           25'b0010011000100010011000100,
           25'b0010001000100010010001000,
           25'b0101001000100010001010100,
           25'b0100001000000000001000100,
           25'b0011001000011100001011000,
           25'b0100001100100010001000100,
           25'b0010000100000000001001000,
           25'b0001100110000000010110000,
           25'b0000011110000001111000000,
           25'b0000000001000010000000000,
           25'b0000000001000100000000000,
           25'b0000000001000100000000000,
           25'b0000000001000100000000000,
           25'b0000000010011000000000000,
           25'b0000000011100000000000000,
           25'b0000000010000000000000000,
           25'b0000000000000000000000000};
    
endmodule 
